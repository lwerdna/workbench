Example from allaboutcircuits.com
v1 1 0 dc 15
r1 1 0 2.2k
r2 1 2 3.3k     
r3 2 0 150
.dc v1 0 15 0.5
.end
